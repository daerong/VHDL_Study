library verilog;
use verilog.vl_types.all;
entity xnor_gate_vlg_vec_tst is
end xnor_gate_vlg_vec_tst;
