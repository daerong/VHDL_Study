library verilog;
use verilog.vl_types.all;
entity MUX_2x1_vlg_vec_tst is
end MUX_2x1_vlg_vec_tst;
