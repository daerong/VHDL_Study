library verilog;
use verilog.vl_types.all;
entity MUX_2x2_vlg_check_tst is
    port(
        Y0              : in     vl_logic;
        Y1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MUX_2x2_vlg_check_tst;
