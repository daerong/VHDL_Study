library verilog;
use verilog.vl_types.all;
entity xor_gate_vlg_vec_tst is
end xor_gate_vlg_vec_tst;
