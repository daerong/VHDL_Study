library verilog;
use verilog.vl_types.all;
entity counter_12_vlg_vec_tst is
end counter_12_vlg_vec_tst;
