library verilog;
use verilog.vl_types.all;
entity FND_Decorder_vlg_vec_tst is
end FND_Decorder_vlg_vec_tst;
