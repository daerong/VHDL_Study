library verilog;
use verilog.vl_types.all;
entity fnd_decoder_vlg_vec_tst is
end fnd_decoder_vlg_vec_tst;
