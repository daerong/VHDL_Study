library verilog;
use verilog.vl_types.all;
entity not_gate_vlg_vec_tst is
end not_gate_vlg_vec_tst;
