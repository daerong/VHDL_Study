library verilog;
use verilog.vl_types.all;
entity MUX_2x1_vlg_check_tst is
    port(
        Y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MUX_2x1_vlg_check_tst;
