library verilog;
use verilog.vl_types.all;
entity xor_gate_vlg_check_tst is
    port(
        pin_name3       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end xor_gate_vlg_check_tst;
