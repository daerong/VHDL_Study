library verilog;
use verilog.vl_types.all;
entity MUX_2x2_vlg_check_tst is
    port(
        Y               : in     vl_logic_vector(1 downto 0);
        sampler_rx      : in     vl_logic
    );
end MUX_2x2_vlg_check_tst;
