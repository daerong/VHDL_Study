library verilog;
use verilog.vl_types.all;
entity DEMUX_1x2_vlg_vec_tst is
end DEMUX_1x2_vlg_vec_tst;
