library verilog;
use verilog.vl_types.all;
entity nand_gate_vlg_vec_tst is
end nand_gate_vlg_vec_tst;
