library verilog;
use verilog.vl_types.all;
entity counter_60_vlg_vec_tst is
end counter_60_vlg_vec_tst;
