library verilog;
use verilog.vl_types.all;
entity MUX_2x2_vlg_vec_tst is
end MUX_2x2_vlg_vec_tst;
