library verilog;
use verilog.vl_types.all;
entity not_gate_vlg_check_tst is
    port(
        pin_name2       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end not_gate_vlg_check_tst;
