library verilog;
use verilog.vl_types.all;
entity nor_gate_vlg_check_tst is
    port(
        Y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end nor_gate_vlg_check_tst;
