library verilog;
use verilog.vl_types.all;
entity DEMUX_1x2_vlg_sample_tst is
    port(
        A               : in     vl_logic;
        SEL             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end DEMUX_1x2_vlg_sample_tst;
