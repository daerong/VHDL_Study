library verilog;
use verilog.vl_types.all;
entity nor_gate_vlg_vec_tst is
end nor_gate_vlg_vec_tst;
